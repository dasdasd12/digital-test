// Copyright (c) 2012 Ben Reynwar
// Released under MIT License (see LICENSE.txt)

module twiddlefactors (
    input  wire                            clk,
    input  wire [7:0]          addr,
    input  wire                            addr_nd,
    output reg signed [19:0] tf_out
  );

  always @ (posedge clk)
    begin
      if (addr_nd)
        begin
          case (addr)
			
            8'd0: tf_out <= { 10'sd256,  -10'sd0 };
			
            8'd1: tf_out <= { 10'sd256,  -10'sd3 };
			
            8'd2: tf_out <= { 10'sd256,  -10'sd6 };
			
            8'd3: tf_out <= { 10'sd256,  -10'sd9 };
			
            8'd4: tf_out <= { 10'sd256,  -10'sd13 };
			
            8'd5: tf_out <= { 10'sd256,  -10'sd16 };
			
            8'd6: tf_out <= { 10'sd255,  -10'sd19 };
			
            8'd7: tf_out <= { 10'sd255,  -10'sd22 };
			
            8'd8: tf_out <= { 10'sd255,  -10'sd25 };
			
            8'd9: tf_out <= { 10'sd254,  -10'sd28 };
			
            8'd10: tf_out <= { 10'sd254,  -10'sd31 };
			
            8'd11: tf_out <= { 10'sd254,  -10'sd34 };
			
            8'd12: tf_out <= { 10'sd253,  -10'sd38 };
			
            8'd13: tf_out <= { 10'sd253,  -10'sd41 };
			
            8'd14: tf_out <= { 10'sd252,  -10'sd44 };
			
            8'd15: tf_out <= { 10'sd252,  -10'sd47 };
			
            8'd16: tf_out <= { 10'sd251,  -10'sd50 };
			
            8'd17: tf_out <= { 10'sd250,  -10'sd53 };
			
            8'd18: tf_out <= { 10'sd250,  -10'sd56 };
			
            8'd19: tf_out <= { 10'sd249,  -10'sd59 };
			
            8'd20: tf_out <= { 10'sd248,  -10'sd62 };
			
            8'd21: tf_out <= { 10'sd248,  -10'sd65 };
			
            8'd22: tf_out <= { 10'sd247,  -10'sd68 };
			
            8'd23: tf_out <= { 10'sd246,  -10'sd71 };
			
            8'd24: tf_out <= { 10'sd245,  -10'sd74 };
			
            8'd25: tf_out <= { 10'sd244,  -10'sd77 };
			
            8'd26: tf_out <= { 10'sd243,  -10'sd80 };
			
            8'd27: tf_out <= { 10'sd242,  -10'sd83 };
			
            8'd28: tf_out <= { 10'sd241,  -10'sd86 };
			
            8'd29: tf_out <= { 10'sd240,  -10'sd89 };
			
            8'd30: tf_out <= { 10'sd239,  -10'sd92 };
			
            8'd31: tf_out <= { 10'sd238,  -10'sd95 };
			
            8'd32: tf_out <= { 10'sd237,  -10'sd98 };
			
            8'd33: tf_out <= { 10'sd235,  -10'sd101 };
			
            8'd34: tf_out <= { 10'sd234,  -10'sd104 };
			
            8'd35: tf_out <= { 10'sd233,  -10'sd107 };
			
            8'd36: tf_out <= { 10'sd231,  -10'sd109 };
			
            8'd37: tf_out <= { 10'sd230,  -10'sd112 };
			
            8'd38: tf_out <= { 10'sd229,  -10'sd115 };
			
            8'd39: tf_out <= { 10'sd227,  -10'sd118 };
			
            8'd40: tf_out <= { 10'sd226,  -10'sd121 };
			
            8'd41: tf_out <= { 10'sd224,  -10'sd123 };
			
            8'd42: tf_out <= { 10'sd223,  -10'sd126 };
			
            8'd43: tf_out <= { 10'sd221,  -10'sd129 };
			
            8'd44: tf_out <= { 10'sd220,  -10'sd132 };
			
            8'd45: tf_out <= { 10'sd218,  -10'sd134 };
			
            8'd46: tf_out <= { 10'sd216,  -10'sd137 };
			
            8'd47: tf_out <= { 10'sd215,  -10'sd140 };
			
            8'd48: tf_out <= { 10'sd213,  -10'sd142 };
			
            8'd49: tf_out <= { 10'sd211,  -10'sd145 };
			
            8'd50: tf_out <= { 10'sd209,  -10'sd147 };
			
            8'd51: tf_out <= { 10'sd207,  -10'sd150 };
			
            8'd52: tf_out <= { 10'sd206,  -10'sd152 };
			
            8'd53: tf_out <= { 10'sd204,  -10'sd155 };
			
            8'd54: tf_out <= { 10'sd202,  -10'sd157 };
			
            8'd55: tf_out <= { 10'sd200,  -10'sd160 };
			
            8'd56: tf_out <= { 10'sd198,  -10'sd162 };
			
            8'd57: tf_out <= { 10'sd196,  -10'sd165 };
			
            8'd58: tf_out <= { 10'sd194,  -10'sd167 };
			
            8'd59: tf_out <= { 10'sd192,  -10'sd170 };
			
            8'd60: tf_out <= { 10'sd190,  -10'sd172 };
			
            8'd61: tf_out <= { 10'sd188,  -10'sd174 };
			
            8'd62: tf_out <= { 10'sd185,  -10'sd177 };
			
            8'd63: tf_out <= { 10'sd183,  -10'sd179 };
			
            8'd64: tf_out <= { 10'sd181,  -10'sd181 };
			
            8'd65: tf_out <= { 10'sd179,  -10'sd183 };
			
            8'd66: tf_out <= { 10'sd177,  -10'sd185 };
			
            8'd67: tf_out <= { 10'sd174,  -10'sd188 };
			
            8'd68: tf_out <= { 10'sd172,  -10'sd190 };
			
            8'd69: tf_out <= { 10'sd170,  -10'sd192 };
			
            8'd70: tf_out <= { 10'sd167,  -10'sd194 };
			
            8'd71: tf_out <= { 10'sd165,  -10'sd196 };
			
            8'd72: tf_out <= { 10'sd162,  -10'sd198 };
			
            8'd73: tf_out <= { 10'sd160,  -10'sd200 };
			
            8'd74: tf_out <= { 10'sd157,  -10'sd202 };
			
            8'd75: tf_out <= { 10'sd155,  -10'sd204 };
			
            8'd76: tf_out <= { 10'sd152,  -10'sd206 };
			
            8'd77: tf_out <= { 10'sd150,  -10'sd207 };
			
            8'd78: tf_out <= { 10'sd147,  -10'sd209 };
			
            8'd79: tf_out <= { 10'sd145,  -10'sd211 };
			
            8'd80: tf_out <= { 10'sd142,  -10'sd213 };
			
            8'd81: tf_out <= { 10'sd140,  -10'sd215 };
			
            8'd82: tf_out <= { 10'sd137,  -10'sd216 };
			
            8'd83: tf_out <= { 10'sd134,  -10'sd218 };
			
            8'd84: tf_out <= { 10'sd132,  -10'sd220 };
			
            8'd85: tf_out <= { 10'sd129,  -10'sd221 };
			
            8'd86: tf_out <= { 10'sd126,  -10'sd223 };
			
            8'd87: tf_out <= { 10'sd123,  -10'sd224 };
			
            8'd88: tf_out <= { 10'sd121,  -10'sd226 };
			
            8'd89: tf_out <= { 10'sd118,  -10'sd227 };
			
            8'd90: tf_out <= { 10'sd115,  -10'sd229 };
			
            8'd91: tf_out <= { 10'sd112,  -10'sd230 };
			
            8'd92: tf_out <= { 10'sd109,  -10'sd231 };
			
            8'd93: tf_out <= { 10'sd107,  -10'sd233 };
			
            8'd94: tf_out <= { 10'sd104,  -10'sd234 };
			
            8'd95: tf_out <= { 10'sd101,  -10'sd235 };
			
            8'd96: tf_out <= { 10'sd98,  -10'sd237 };
			
            8'd97: tf_out <= { 10'sd95,  -10'sd238 };
			
            8'd98: tf_out <= { 10'sd92,  -10'sd239 };
			
            8'd99: tf_out <= { 10'sd89,  -10'sd240 };
			
            8'd100: tf_out <= { 10'sd86,  -10'sd241 };
			
            8'd101: tf_out <= { 10'sd83,  -10'sd242 };
			
            8'd102: tf_out <= { 10'sd80,  -10'sd243 };
			
            8'd103: tf_out <= { 10'sd77,  -10'sd244 };
			
            8'd104: tf_out <= { 10'sd74,  -10'sd245 };
			
            8'd105: tf_out <= { 10'sd71,  -10'sd246 };
			
            8'd106: tf_out <= { 10'sd68,  -10'sd247 };
			
            8'd107: tf_out <= { 10'sd65,  -10'sd248 };
			
            8'd108: tf_out <= { 10'sd62,  -10'sd248 };
			
            8'd109: tf_out <= { 10'sd59,  -10'sd249 };
			
            8'd110: tf_out <= { 10'sd56,  -10'sd250 };
			
            8'd111: tf_out <= { 10'sd53,  -10'sd250 };
			
            8'd112: tf_out <= { 10'sd50,  -10'sd251 };
			
            8'd113: tf_out <= { 10'sd47,  -10'sd252 };
			
            8'd114: tf_out <= { 10'sd44,  -10'sd252 };
			
            8'd115: tf_out <= { 10'sd41,  -10'sd253 };
			
            8'd116: tf_out <= { 10'sd38,  -10'sd253 };
			
            8'd117: tf_out <= { 10'sd34,  -10'sd254 };
			
            8'd118: tf_out <= { 10'sd31,  -10'sd254 };
			
            8'd119: tf_out <= { 10'sd28,  -10'sd254 };
			
            8'd120: tf_out <= { 10'sd25,  -10'sd255 };
			
            8'd121: tf_out <= { 10'sd22,  -10'sd255 };
			
            8'd122: tf_out <= { 10'sd19,  -10'sd255 };
			
            8'd123: tf_out <= { 10'sd16,  -10'sd256 };
			
            8'd124: tf_out <= { 10'sd13,  -10'sd256 };
			
            8'd125: tf_out <= { 10'sd9,  -10'sd256 };
			
            8'd126: tf_out <= { 10'sd6,  -10'sd256 };
			
            8'd127: tf_out <= { 10'sd3,  -10'sd256 };
			
            8'd128: tf_out <= { 10'sd0,  -10'sd256 };
			
            8'd129: tf_out <= { -10'sd3,  -10'sd256 };
			
            8'd130: tf_out <= { -10'sd6,  -10'sd256 };
			
            8'd131: tf_out <= { -10'sd9,  -10'sd256 };
			
            8'd132: tf_out <= { -10'sd13,  -10'sd256 };
			
            8'd133: tf_out <= { -10'sd16,  -10'sd256 };
			
            8'd134: tf_out <= { -10'sd19,  -10'sd255 };
			
            8'd135: tf_out <= { -10'sd22,  -10'sd255 };
			
            8'd136: tf_out <= { -10'sd25,  -10'sd255 };
			
            8'd137: tf_out <= { -10'sd28,  -10'sd254 };
			
            8'd138: tf_out <= { -10'sd31,  -10'sd254 };
			
            8'd139: tf_out <= { -10'sd34,  -10'sd254 };
			
            8'd140: tf_out <= { -10'sd38,  -10'sd253 };
			
            8'd141: tf_out <= { -10'sd41,  -10'sd253 };
			
            8'd142: tf_out <= { -10'sd44,  -10'sd252 };
			
            8'd143: tf_out <= { -10'sd47,  -10'sd252 };
			
            8'd144: tf_out <= { -10'sd50,  -10'sd251 };
			
            8'd145: tf_out <= { -10'sd53,  -10'sd250 };
			
            8'd146: tf_out <= { -10'sd56,  -10'sd250 };
			
            8'd147: tf_out <= { -10'sd59,  -10'sd249 };
			
            8'd148: tf_out <= { -10'sd62,  -10'sd248 };
			
            8'd149: tf_out <= { -10'sd65,  -10'sd248 };
			
            8'd150: tf_out <= { -10'sd68,  -10'sd247 };
			
            8'd151: tf_out <= { -10'sd71,  -10'sd246 };
			
            8'd152: tf_out <= { -10'sd74,  -10'sd245 };
			
            8'd153: tf_out <= { -10'sd77,  -10'sd244 };
			
            8'd154: tf_out <= { -10'sd80,  -10'sd243 };
			
            8'd155: tf_out <= { -10'sd83,  -10'sd242 };
			
            8'd156: tf_out <= { -10'sd86,  -10'sd241 };
			
            8'd157: tf_out <= { -10'sd89,  -10'sd240 };
			
            8'd158: tf_out <= { -10'sd92,  -10'sd239 };
			
            8'd159: tf_out <= { -10'sd95,  -10'sd238 };
			
            8'd160: tf_out <= { -10'sd98,  -10'sd237 };
			
            8'd161: tf_out <= { -10'sd101,  -10'sd235 };
			
            8'd162: tf_out <= { -10'sd104,  -10'sd234 };
			
            8'd163: tf_out <= { -10'sd107,  -10'sd233 };
			
            8'd164: tf_out <= { -10'sd109,  -10'sd231 };
			
            8'd165: tf_out <= { -10'sd112,  -10'sd230 };
			
            8'd166: tf_out <= { -10'sd115,  -10'sd229 };
			
            8'd167: tf_out <= { -10'sd118,  -10'sd227 };
			
            8'd168: tf_out <= { -10'sd121,  -10'sd226 };
			
            8'd169: tf_out <= { -10'sd123,  -10'sd224 };
			
            8'd170: tf_out <= { -10'sd126,  -10'sd223 };
			
            8'd171: tf_out <= { -10'sd129,  -10'sd221 };
			
            8'd172: tf_out <= { -10'sd132,  -10'sd220 };
			
            8'd173: tf_out <= { -10'sd134,  -10'sd218 };
			
            8'd174: tf_out <= { -10'sd137,  -10'sd216 };
			
            8'd175: tf_out <= { -10'sd140,  -10'sd215 };
			
            8'd176: tf_out <= { -10'sd142,  -10'sd213 };
			
            8'd177: tf_out <= { -10'sd145,  -10'sd211 };
			
            8'd178: tf_out <= { -10'sd147,  -10'sd209 };
			
            8'd179: tf_out <= { -10'sd150,  -10'sd207 };
			
            8'd180: tf_out <= { -10'sd152,  -10'sd206 };
			
            8'd181: tf_out <= { -10'sd155,  -10'sd204 };
			
            8'd182: tf_out <= { -10'sd157,  -10'sd202 };
			
            8'd183: tf_out <= { -10'sd160,  -10'sd200 };
			
            8'd184: tf_out <= { -10'sd162,  -10'sd198 };
			
            8'd185: tf_out <= { -10'sd165,  -10'sd196 };
			
            8'd186: tf_out <= { -10'sd167,  -10'sd194 };
			
            8'd187: tf_out <= { -10'sd170,  -10'sd192 };
			
            8'd188: tf_out <= { -10'sd172,  -10'sd190 };
			
            8'd189: tf_out <= { -10'sd174,  -10'sd188 };
			
            8'd190: tf_out <= { -10'sd177,  -10'sd185 };
			
            8'd191: tf_out <= { -10'sd179,  -10'sd183 };
			
            8'd192: tf_out <= { -10'sd181,  -10'sd181 };
			
            8'd193: tf_out <= { -10'sd183,  -10'sd179 };
			
            8'd194: tf_out <= { -10'sd185,  -10'sd177 };
			
            8'd195: tf_out <= { -10'sd188,  -10'sd174 };
			
            8'd196: tf_out <= { -10'sd190,  -10'sd172 };
			
            8'd197: tf_out <= { -10'sd192,  -10'sd170 };
			
            8'd198: tf_out <= { -10'sd194,  -10'sd167 };
			
            8'd199: tf_out <= { -10'sd196,  -10'sd165 };
			
            8'd200: tf_out <= { -10'sd198,  -10'sd162 };
			
            8'd201: tf_out <= { -10'sd200,  -10'sd160 };
			
            8'd202: tf_out <= { -10'sd202,  -10'sd157 };
			
            8'd203: tf_out <= { -10'sd204,  -10'sd155 };
			
            8'd204: tf_out <= { -10'sd206,  -10'sd152 };
			
            8'd205: tf_out <= { -10'sd207,  -10'sd150 };
			
            8'd206: tf_out <= { -10'sd209,  -10'sd147 };
			
            8'd207: tf_out <= { -10'sd211,  -10'sd145 };
			
            8'd208: tf_out <= { -10'sd213,  -10'sd142 };
			
            8'd209: tf_out <= { -10'sd215,  -10'sd140 };
			
            8'd210: tf_out <= { -10'sd216,  -10'sd137 };
			
            8'd211: tf_out <= { -10'sd218,  -10'sd134 };
			
            8'd212: tf_out <= { -10'sd220,  -10'sd132 };
			
            8'd213: tf_out <= { -10'sd221,  -10'sd129 };
			
            8'd214: tf_out <= { -10'sd223,  -10'sd126 };
			
            8'd215: tf_out <= { -10'sd224,  -10'sd123 };
			
            8'd216: tf_out <= { -10'sd226,  -10'sd121 };
			
            8'd217: tf_out <= { -10'sd227,  -10'sd118 };
			
            8'd218: tf_out <= { -10'sd229,  -10'sd115 };
			
            8'd219: tf_out <= { -10'sd230,  -10'sd112 };
			
            8'd220: tf_out <= { -10'sd231,  -10'sd109 };
			
            8'd221: tf_out <= { -10'sd233,  -10'sd107 };
			
            8'd222: tf_out <= { -10'sd234,  -10'sd104 };
			
            8'd223: tf_out <= { -10'sd235,  -10'sd101 };
			
            8'd224: tf_out <= { -10'sd237,  -10'sd98 };
			
            8'd225: tf_out <= { -10'sd238,  -10'sd95 };
			
            8'd226: tf_out <= { -10'sd239,  -10'sd92 };
			
            8'd227: tf_out <= { -10'sd240,  -10'sd89 };
			
            8'd228: tf_out <= { -10'sd241,  -10'sd86 };
			
            8'd229: tf_out <= { -10'sd242,  -10'sd83 };
			
            8'd230: tf_out <= { -10'sd243,  -10'sd80 };
			
            8'd231: tf_out <= { -10'sd244,  -10'sd77 };
			
            8'd232: tf_out <= { -10'sd245,  -10'sd74 };
			
            8'd233: tf_out <= { -10'sd246,  -10'sd71 };
			
            8'd234: tf_out <= { -10'sd247,  -10'sd68 };
			
            8'd235: tf_out <= { -10'sd248,  -10'sd65 };
			
            8'd236: tf_out <= { -10'sd248,  -10'sd62 };
			
            8'd237: tf_out <= { -10'sd249,  -10'sd59 };
			
            8'd238: tf_out <= { -10'sd250,  -10'sd56 };
			
            8'd239: tf_out <= { -10'sd250,  -10'sd53 };
			
            8'd240: tf_out <= { -10'sd251,  -10'sd50 };
			
            8'd241: tf_out <= { -10'sd252,  -10'sd47 };
			
            8'd242: tf_out <= { -10'sd252,  -10'sd44 };
			
            8'd243: tf_out <= { -10'sd253,  -10'sd41 };
			
            8'd244: tf_out <= { -10'sd253,  -10'sd38 };
			
            8'd245: tf_out <= { -10'sd254,  -10'sd34 };
			
            8'd246: tf_out <= { -10'sd254,  -10'sd31 };
			
            8'd247: tf_out <= { -10'sd254,  -10'sd28 };
			
            8'd248: tf_out <= { -10'sd255,  -10'sd25 };
			
            8'd249: tf_out <= { -10'sd255,  -10'sd22 };
			
            8'd250: tf_out <= { -10'sd255,  -10'sd19 };
			
            8'd251: tf_out <= { -10'sd256,  -10'sd16 };
			
            8'd252: tf_out <= { -10'sd256,  -10'sd13 };
			
            8'd253: tf_out <= { -10'sd256,  -10'sd9 };
			
            8'd254: tf_out <= { -10'sd256,  -10'sd6 };
			
            8'd255: tf_out <= { -10'sd256,  -10'sd3 };
			
            default:
              begin
                tf_out <= 20'd0;
              end
         endcase
      end
  end
endmodule